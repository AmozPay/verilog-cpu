
module tb_dmux;
endmodule