
module tb_or_nway;
endmodule