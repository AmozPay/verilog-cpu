`include "src/boolean/xor_nbits.v"
// Perfom xor between two buses
module tb_xor_nbits;
endmodule
