`include "src/boolean/and_nway.v"

module tb_nand_nbits;
endmodule
