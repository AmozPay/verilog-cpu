
// Perfom or between two buses
module tb_or_nbits;

endmodule