`include "src/boolean/and_nway.v"

module tb_and_nbits;
endmodule
